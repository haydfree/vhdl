library IEEE;
use IEEE.std_logic_1164.all;

entity tb is
end entity;

architecture test of tb is

begin

end architecture;

library IEEE;
use IEEE.std_logic_1164.all;

entity HACK_NOT is

end entity;

architecture rtl of HACK_NOT is

begin

end architecture;
